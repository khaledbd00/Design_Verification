module counter(
	input [15:0] data_in,
	input clk,
	input reset,
	input load,
	input enable,
	input up_down,
	output [15:0] data_out
	);
endmodule